module pc_sel (
    input wire Zero, Gt, PCWrite, PCWriteCond, EQorNE, GTorLT,
    output wire Out
);

    wire notZero, notGt;
    wire rZeroGt, rAux;
	 wire EQorNE_Out, GTorLT_Out;
	 

    assign notZero = ~Zero;
    assign notGt = ~Gt;

    mux_2x1_1_1 Mux_EQorNE(EQorNE_Out, EQorNE, notZero, Zero); 
    mux_2x1_1_1 Mux_GTorLT(GTorLT_Out, GTorLT, notGt, Gt); 
	 

    assign rZeroGt = EQorNE_Out | GTorLT_Out;
    assign rAux = rZeroGt & PCWriteCond;
    assign Out = rAux | PCWrite;
    
endmodule