module controladora (
    ports
);
    
endmodule